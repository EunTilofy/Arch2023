`timescale 1ns / 1ps

module core_sim;
    reg clk, rst;

    initial begin
        $dumpfile("wave.vcd");
        $dumpvars;
        #1000
        $finish;
    end

    RV32core core(
        .debug_en(1'b0),
        .debug_step(1'b0),
        .debug_addr(7'b0),
        .debug_data(),
        .clk(clk),
        .rst(rst),
        .interrupter(1'b0)
    );

    initial begin
        clk = 0;
        rst = 1;
        #2 rst = 0;
    end
    always #1 clk = ~clk;

endmodule